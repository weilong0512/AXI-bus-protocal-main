`include "SRAM.sv"

