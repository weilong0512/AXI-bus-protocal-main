`define DATAWIDTH 32 
`define SIZE 3 